`include "test_scenario_base.sv"

`include "axi_rw_000.sv"
